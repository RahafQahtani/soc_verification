
`define SPI1_BASE_ADDRESS 32'h20000200
`define SPI1_END_ADDRESS 32'h2000027F
`define SPI2_BASE_ADDRESS 32'h20000280
`define SPI2_END_ADDRESS 32'h200002FF
`define OFFSET 4
